library ieee;
use ieee.std_logic_1164.all;

entity blub is
port(
      TX_DATA  : out std_logic_vector(1 downto 0) --TODO

);
end entity blub;
