test file
blub
blubblub
