library ieee;
use ieee.std_logic_1164.all;

entity blub is
port(


);
end entity blub;
