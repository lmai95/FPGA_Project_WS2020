test file
blub
blub2
